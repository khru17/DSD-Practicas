LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY palabra IS PORT (
    CLR, CLK, EN : IN STD_LOGIC;
    DISPLAY : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
ATTRIBUTE PIN_NUMBERS OF palabra : ENTITY IS
"CLK:1 EN:2 CLR:13 DISPLAY(6):23 DISPLAY(5):22 DISPLAY(4):21 DISPLAY(3):20 DISPLAY(2):19 DISPLAY(1):18 DISPLAY(0):17";
END palabra;

ARCHITECTURE A_palabra OF palabra IS
-- ALIAS
CONSTANT L0 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
CONSTANT L1 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
CONSTANT L2 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
-- LETRAS
CONSTANT H : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110111";
CONSTANT O : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1111110";
CONSTANT L : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001110";
CONSTANT A : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110111";
CONSTANT S : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1011011";
CONSTANT I : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
CONSTANT G : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1011111";
CONSTANT C : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001110";
CONSTANT U : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0111110";
CONSTANT B : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0011111";
-- SE�AL DE APOYO
SIGNAL SAL : STD_LOGIC_VECTOR(8 DOWNTO 0);
-- LETRA CON SU ALIAS
CONSTANT EH_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&H;
CONSTANT EO_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&O;
CONSTANT EL_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&L;
CONSTANT EA_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&A;
CONSTANT ES_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&S;
CONSTANT EO_1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L1&O;
CONSTANT EI_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&I;
CONSTANT EG_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&G;
CONSTANT EO_2 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L2&O;
CONSTANT EC_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&C;
CONSTANT EU_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&U;
CONSTANT EB_0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L0&B;
CONSTANT EA_1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L1&A;
CONSTANT EI_1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := L1&I;

BEGIN
    PROCESS (CLK, CLR)
    BEGIN
        IF (CLR = '1') THEN
            SAL <= EH_0;
        ELSIF ( RISING_EDGE(CLK)) THEN
            IF ( EN = '1' ) THEN
                CASE SAL IS 
                    WHEN EH_0 => SAL <= EO_0;
                    WHEN EO_0 => SAL <= EL_0;
                    WHEN EL_0 => SAL <= EA_0;
                    WHEN EA_0 => SAL <= ES_0;
                    WHEN ES_0 => SAL <= EO_1;
                    WHEN EO_1 => SAL <= EI_0;
                    WHEN EI_0 => SAL <= EG_0;
                    WHEN EG_0 => SAL <= EO_2;
                    WHEN EO_2 => SAL <= EC_0;
                    WHEN EC_0 => SAL <= EU_0;
                    WHEN EU_0 => SAL <= EB_0;
                    WHEN EB_0 => SAL <= EA_1;
                    WHEN EA_1 => SAL <= EI_1;
                    WHEN EI_1 => SAL <= EH_0;
                    WHEN OTHERS => SAL <= EH_0;
                END CASE;
            END IF;
        END IF;
    END PROCESS;

    DISPLAY <= SAL(6 DOWNTO 0);

END A_palabra;