module multiplexer ( 
	clk,
	clr,
	display,
	sel
	) ;

input  clk;
input  clr;
inout [6:0] display;
inout [2:0] sel;
