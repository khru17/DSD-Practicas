module p2 ( 
	d,
	t,
	s,
	r,
	j,
	k,
	clk,
	clr,
	sel,
	sal
	) ;

input  d;
input  t;
input  s;
input  r;
input  j;
input  k;
input  clk;
input  clr;
input [1:0] sel;
inout [5:0] sal;
