LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY teclado IS PORT (
    CLR, CLK, L : IN STD_LOGIC;
    DISPLAY : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    COLUMNA : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    FILA: IN STD_LOGIC_VECTOR(3 DOWNTO 0)
);
ATTRIBUTE PIN_NUMBERS OF teclado : ENTITY IS
    "CLK:1 L:2 FILA(3):5 FILA(2):6 FILA(1):7 FILA(0):8, CLR:13 "&
    "COLUMNA(2):23 COLUMNA(1):22 COLUMNA(0):21 "&
    "DISPLAY(6):20 DISPLAY(5):19 DISPLAY(4):18 DISPLAY(3):17 DISPLAY(2):16 "&
    "DISPLAY(1):15 DISPLAY(0):14";
END teclado;

ARCHITECTURE A_teclado OF teclado IS

CONSTANT N0 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1111110"; -- 7E
CONSTANT N1 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "0110000"; -- 30
CONSTANT N2 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1101101"; -- 6D
CONSTANT N3 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1111001"; -- 79
CONSTANT N4 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "0110011"; -- 33
CONSTANT N5 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1011011"; -- 5B
CONSTANT N6 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "0011111"; -- 1F
CONSTANT N7 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1110000"; -- 70
CONSTANT N8 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1111111"; -- 7F
CONSTANT N9 : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1110011"; -- 73
CONSTANT N_A : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "1110111"; -- 77
CONSTANT N_H : STD_LOGIC_VECTOR (6 DOWNTO 0 ) := "0110111"; -- 37

SIGNAL D: STD_LOGIC_VECTOR(6 DOWNTO 0);

BEGIN
    -- CONTADOR DE ANILLO CON 0 VIAJERO
    ANILLO : PROCESS ( CLR, CLK )
    BEGIN
        IF ( CLR = '1' ) THEN
            COLUMNA <= "011";
        ELSIF ( CLK'EVENT AND CLK = '1' ) THEN  
            CASE COLUMNA IS
				WHEN "011" => COLUMNA <= "101";
				WHEN "101" => COLUMNA <= "110";
				WHEN "110" => COLUMNA <= "011";
				WHEN OTHERS => COLUMNA <= "---";
			END CASE;
        END IF;
    END PROCESS ANILLO;

    -- DECODIFICADOR
    DECODIFICADOR : PROCESS ( COLUMNA, FILA )
    BEGIN
        CASE FILA&COLUMNA IS
            WHEN "1110011" => D <= N1;
            WHEN "1110101" => D <= N2;
            WHEN "1110110" => D <= N3;

            WHEN "1101011" => D <= N4;
            WHEN "1101101" => D <= N5;
            WHEN "1101110" => D <= N6;

            WHEN "1011011" => D <= N7;
            WHEN "1011101" => D <= N8;
            WHEN "1011110" => D <= N9;

            WHEN "0111011" => D <= N_A;
            WHEN "0111101" => D <= N0;
            WHEN "0111110" => D <= N_H;
            WHEN OTHERS => D <= "-------";
        END CASE;
    END PROCESS DECODIFICADOR;

    -- REGISTRO
    REGISTRO : PROCESS ( CLR, CLK )
    BEGIN
        IF ( CLR = '1' ) THEN
            DISPLAY<=(OTHERS=>'0');
        ELSIF ( CLK'EVENT AND CLK = '1' ) THEN 
            IF(L='1') THEN  
                DISPLAY <= D;
            ELSE    
                DISPLAY <= DISPLAY;
            END IF;
        END IF;
    END PROCESS REGISTRO;

END A_teclado;