module p3 ( 
	d,
	es,
	clk,
	clr,
	sel,
	q
	) ;

input [6:0] d;
input  es;
input  clk;
input  clr;
input [1:0] sel;
inout [6:0] q;
