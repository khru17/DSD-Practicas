module contador ( 
	en,
	clk,
	clr,
	q
	) ;

input  en;
input  clk;
input  clr;
inout [2:0] q;
