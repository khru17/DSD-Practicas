module palabra ( 
	clr,
	clk,
	en,
	display
	) ;

input  clr;
input  clk;
input  en;
inout [6:0] display;
