module practica1 ( 
	a,
	b,
	ref,
	sel,
	comparador,
	display
	) ;

input [2:0] a;
input [2:0] b;
input [2:0] ref;
input  sel;
inout [2:0] comparador;
inout [6:0] display;
