module sensores_1 ( 
	unid,
	dece,
	ent,
	clr,
	clk
	) ;

inout [3:0] unid;
inout [2:0] dece;
input [1:0] ent;
input  clr;
input  clk;
