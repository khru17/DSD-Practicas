module sensores_2 ( 
	clr,
	clk,
	display,
	unid,
	dece,
	sel
	) ;

input  clr;
input  clk;
inout [6:0] display;
input [3:0] unid;
input [2:0] dece;
inout [2:0] sel;
