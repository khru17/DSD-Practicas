module cartaasm ( 
	d,
	clk,
	clr,
	ini,
	a,
	lb,
	eb,
	ec
	) ;

input [5:0] d;
input  clk;
input  clr;
input  ini;
inout [5:0] a;
inout  lb;
inout  eb;
inout  ec;
