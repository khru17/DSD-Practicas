module mealy ( 
	clk,
	clr,
	e,
	sal,
	display
	) ;

input  clk;
input  clr;
input  e;
inout  sal;
inout [6:0] display;
