module contador_10 ( 
	clk,
	clr,
	e,
	q
	) ;

input  clk;
input  clr;
input  e;
inout [9:0] q;
